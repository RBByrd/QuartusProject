LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY main IS 
PORT(
 clock, reset : IN STD_LOGIC; 
 IR2o : OUT STD_LOGIC_VECTOR(31 DOWNTO 0 ); 
 PC2o  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0 );
 IR3o : OUT STD_LOGIC_VECTOR (13 DOWNTO 0); 
 X3o  : out STD_LOGIC_VECTOR (31 DOWNTO 0);    
 Y3o  : OUT STD_LOGIC_VECTOR (31 DOWNTO 0); 
 MD3o  : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
 IR4o : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);     
 Z4o  : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
 MD4o  : out STD_LOGIC_VECTOR (31 DOWNTO 0);
 IR5o : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);  
 MP1o  : OUT STD_LOGIC;
 Z5o  : out STD_LOGIC_VECTOR (31 DOWNTO 0) 
 	
);
end main;

ARCHITECTURE a OF main IS

signal IR2 : STD_LOGIC_VECTOR(31 DOWNTO 0 );
signal PC2  :  STD_LOGIC_VECTOR(31 DOWNTO 0 );
signal 	MP1 :  STD_LOGIC;
signal 	RB :  STD_LOGIC_VECTOR (31 DOWNTO 0);
signal IR3	: STD_LOGIC_VECTOR(13 DOWNTO 0);
signal X3   :  STD_LOGIC_VECTOR(31 DOWNTO 0);
signal 	Y3 :STD_LOGIC_VECTOR(31 DOWNTO 0);
signal 	R1		: STD_LOGIC_VECTOR(31 DOWNTO 0);
signal 	R2		: STD_LOGIC_VECTOR(31 DOWNTO 0);
signal	MP2 :  STD_LOGIC;
signal	MD3 : STD_LOGIC_VECTOR(31 DOWNTO 0);
signal	IR5 	:  STD_LOGIC_VECTOR(7 DOWNTO 0);
signal	Z5		:  STD_LOGIC_VECTOR(31 DOWNTO 0);
signal	w3		:  STD_LOGIC;
signal   MD4 :  STD_LOGIC_VECTOR (31 DOWNTO 0); 
signal	   IR4 :  STD_LOGIC_VECTOR (7 DOWNTO 0); 
signal   Z4 :  STD_LOGIC_VECTOR (31 DOWNTO 0); 
signal MP7 :  STD_LOGIC_VECTOR (1 DOWNTO 0); 
signal MP6 :  STD_LOGIC_VECTOR (1 DOWNTO 0); 
signal	MD3i : STD_LOGIC_VECTOR(31 DOWNTO 0);  

component fetch 
PORT( 
	clock, reset : IN STD_LOGIC; 
	IR2 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0 ); 
	PC2  : OUT STD_LOGIC_VECTOR(31 DOWNTO 0 );
	MP1 : in STD_LOGIC;
	RB : IN STD_LOGIC_VECTOR (31 DOWNTO 0));

   END component;
component vhdl1 --decode
PORT(
	CLOCK : IN STD_LOGIC;
	RESET : IN STD_LOGIC;
	IR2	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	PC2   : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	IR3	: OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
	X3		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	Y3 	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	R1		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	R2		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	MP2 : OUT STD_LOGIC;
	MD3 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	MP1 : OUT STD_LOGIC
	
	);
end component;
	component RF 
PORT(
	CLOCK : IN STD_LOGIC;
	RESET : IN STD_LOGIC;
	IR2	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	IR5 	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	Z5		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	w3		: IN STD_LOGIC;

	R1	   : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	R2		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	MP2 	: IN STD_LOGIC;
	MD3 	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
  end component;	
  component MEM_ACCESS
PORT( 
	clock, reset : IN STD_LOGIC; 
   IR4 : IN STD_LOGIC_VECTOR (7 DOWNTO 0); 
   Z4 : IN STD_LOGIC_VECTOR (31 DOWNTO 0); 
   MD4 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);  
   IR5 : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);	
   Z5  : OUT STD_LOGIC_VECTOR (31 DOWNTO 0) 
   ); 
END component;
component Arithmetic_Logic_Unit      
PORT(     
	clock, reset : IN STD_LOGIC;   
	IR3 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);     
	X3  : IN STD_LOGIC_VECTOR (31 DOWNTO 0);    
	Y3  : IN STD_LOGIC_VECTOR (31 DOWNTO 0);  
	Z5  : IN STD_LOGIC_VECTOR (31 DOWNTO 0);    
	MD3 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);   
	Z4 : IN STD_LOGIC_VECTOR (31 DOWNTO 0);   
	MP6 : IN STD_LOGIC_VECTOR (1 DOWNTO 0);   
	MP7 : IN STD_LOGIC_VECTOR (1 DOWNTO 0);   
	IR4 : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);   
	C : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);   
	MD4 : OUT STD_LOGIC_VECTOR (31 DOWNTO 0)   
  );     
END component;


component RA_WRITE IS
PORT(
	CLOCK : IN STD_LOGIC;
	RESET : IN STD_LOGIC;
	IR5 : IN STD_LOGIC_VECTOR (7 DOWNTO 0);
	Z5 : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
--	A3 : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
--	R3 : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
	W3 : OUT STD_LOGIC
	);
  end component;
	
	component hazards01 IS
PORT(
	CLOCK : IN STD_LOGIC;
	RESET : IN STD_LOGIC;
	IR3 : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
	IR4 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	MPB : OUT STD_LOGIC;
	MPC : OUT STD_LOGIC
	);
  end component;
  
  component hazards02 IS
PORT(
	CLOCK : IN STD_LOGIC;
	RESET : IN STD_LOGIC;
	IR3 : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
	IR5 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	MPB : OUT STD_LOGIC;
	MPC : OUT STD_LOGIC
	);
  end component;
	
	BEGIN
	
		IR2o <= IR2;
		PC2o  <= Pc2;
		IR3o <= IR3;
		X3o  <= X3 ;  
		Y3o  <= Y3 ; 
		MD3o <= MD3i;	
		IR4o <= IR4;    
		Z4o  <= Z4;
		MD4o  <= MD4;
		IR5o <= IR5;    
		Z5o  <= Z5;
		MD3 <= MD3i;
		mp1o <= mp1;		
		
	
		C1 : fetch port map ( Clock ,reset,
		IR2, PC2, MP1, X3);
		C2 : vhdl1 PORT MAP (Clock ,reset,         --decode
		IR2, PC2 , IR3, X3, Y3, R1, R2, MP2, MD3 , MP1);
		C3 : RF PORT MAP(CLOCK, RESET, IR2 , IR5, Z5, w3,
		R1, R2, MP2, MD3);
		C4 : MEM_ACCESS PORT MAP (clock, reset, IR4, Z4,
		MD4, IR5, Z5);
		C5 : Arithmetic_Logic_Unit Port Map (clock, reset, IR3(13 DOWNTO 6), X3, Y3,
		Z5, MD3i, Z4, MP6, MP7, IR4, Z4, MD4);
		C6 : RA_WRITE PORT MAP (Clock, Reset, IR5, Z5, W3);
		C7 : hazards01 PORT MAP (CLock, Reset, IR3(5 downto 0), IR4, MP6(1), MP7(1));
		C8 : hazards02 PORT MAP (CLOCK, RESET, IR3(5 downto 0), IR5, MP6(0), MP7(0));


	
END ARCHITECTURE;
