LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY RF IS
PORT(
	CLOCK : IN STD_LOGIC;
	RESET : IN STD_LOGIC;
	IR2	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	IR5 	: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	Z5		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	w3		: IN STD_LOGIC;

	R1	   : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	R2		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	
	MP2 	: IN STD_LOGIC;
	MD3 	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
  end RF;

 
ARCHITECTURE a OF RF IS 

TYPE reg_file IS array (0 DOWNTO 7) of STD_LOGIC_VECTOR(31 DOWNTO 0);
 SIGNAL R: reg_file;

 
  Begin
	
	PROCESS(CLOCK, RESET)
	begin
		IF reset = '1' THEN
		
			R1(31 DOWNTO 0) <= R(CONV_INTEGER(IR2(21 DOWNTO 19))); --R1
			
			
			--MP2
			CASE MP2 IS
				WHEN '0' => --R[ra]
					R2(31 DOWNTO 0) <= R(CONV_INTEGER(IR2(20 DOWNTO 18))); --rc
			   WHEN '1' => --R[rb]
					R2(31 DOWNTO 0) <= R(CONV_INTEGER(IR2(26 DOWNTO 24))); --ra
				WHEN OTHERS =>
				END CASE;
			
			--W3
			CASE W3 IS 
				WHEN '1' => --load
				R(CONV_INTEGER(IR5(2 DOWNTO 0))) <= Z5; 
			WHEN OTHERS =>
			END CASE;
			end if;	
				
	END PROCESS;
END ARCHITECTURE;